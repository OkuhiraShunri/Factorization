`timescale 1ns / 100ps

module DB_SIM();

reg clk;
reg [3:0] num;
wire [23:0] que;

DB d0(
    .CLK(clk),
    .NUM_IN(num),
    .QUESTION(que)
);

always begin
        clk = 1;
  #0.8  clk = 0;
  #0.8;
end


initial begin
    num = 4'd4;
  #50 num = 4'd0;
end

endmodule